magic
tech sky130A
timestamp 1695672883
<< nwell >>
rect -145 585 280 895
rect -125 535 35 585
rect -125 270 30 535
<< nmos >>
rect -55 -165 -40 235
rect -5 135 10 235
rect 150 420 165 520
rect 150 290 165 390
rect -5 -165 10 -65
rect 190 115 205 215
rect 190 -80 205 20
<< pmos >>
rect -75 775 -60 875
rect 150 775 165 875
rect 190 775 205 875
rect -55 605 -40 705
rect -55 420 -40 520
rect -55 290 -40 390
rect 150 605 165 705
rect 190 605 205 705
<< ndiff >>
rect -105 220 -55 235
rect -105 -150 -90 220
rect -70 -150 -55 220
rect -105 -165 -55 -150
rect -40 135 -5 235
rect 10 220 60 235
rect 10 150 25 220
rect 45 150 60 220
rect 10 135 60 150
rect -40 -65 -15 135
rect 100 505 150 520
rect 100 435 115 505
rect 135 435 150 505
rect 100 420 150 435
rect 165 505 215 520
rect 165 435 180 505
rect 200 435 215 505
rect 165 420 215 435
rect 100 375 150 390
rect 100 305 115 375
rect 135 305 150 375
rect 100 290 150 305
rect 165 375 215 390
rect 165 305 180 375
rect 200 305 215 375
rect 165 290 215 305
rect -40 -165 -5 -65
rect 10 -80 60 -65
rect 10 -150 25 -80
rect 45 -150 60 -80
rect 10 -165 60 -150
rect 140 200 190 215
rect 140 130 155 200
rect 175 130 190 200
rect 140 115 190 130
rect 205 200 255 215
rect 205 130 220 200
rect 240 130 255 200
rect 205 115 255 130
rect 140 5 190 20
rect 140 -65 155 5
rect 175 -65 190 5
rect 140 -80 190 -65
rect 205 5 255 20
rect 205 -65 220 5
rect 240 -65 255 5
rect 205 -80 255 -65
<< pdiff >>
rect -125 860 -75 875
rect -125 790 -110 860
rect -90 790 -75 860
rect -125 775 -75 790
rect -60 860 -10 875
rect -60 790 -45 860
rect -25 790 -10 860
rect -60 775 -10 790
rect 100 860 150 875
rect 100 790 115 860
rect 135 790 150 860
rect 100 775 150 790
rect 165 775 190 875
rect 205 860 255 875
rect 205 790 220 860
rect 240 790 255 860
rect 205 775 255 790
rect -105 690 -55 705
rect -105 620 -90 690
rect -70 620 -55 690
rect -105 605 -55 620
rect -40 690 10 705
rect -40 620 -25 690
rect -5 620 10 690
rect -40 605 10 620
rect -105 505 -55 520
rect -105 435 -90 505
rect -70 435 -55 505
rect -105 420 -55 435
rect -40 505 10 520
rect -40 435 -25 505
rect -5 435 10 505
rect -40 420 10 435
rect -105 375 -55 390
rect -105 305 -90 375
rect -70 305 -55 375
rect -105 290 -55 305
rect -40 375 10 390
rect -40 305 -25 375
rect -5 305 10 375
rect -40 290 10 305
rect 100 690 150 705
rect 100 620 115 690
rect 135 620 150 690
rect 100 605 150 620
rect 165 605 190 705
rect 205 690 255 705
rect 205 620 220 690
rect 240 620 255 690
rect 205 605 255 620
<< ndiffc >>
rect -90 -150 -70 220
rect 25 150 45 220
rect 115 435 135 505
rect 180 435 200 505
rect 115 305 135 375
rect 180 305 200 375
rect 25 -150 45 -80
rect 155 130 175 200
rect 220 130 240 200
rect 155 -65 175 5
rect 220 -65 240 5
<< pdiffc >>
rect -110 790 -90 860
rect -45 790 -25 860
rect 115 790 135 860
rect 220 790 240 860
rect -90 620 -70 690
rect -25 620 -5 690
rect -90 435 -70 505
rect -25 435 -5 505
rect -90 305 -70 375
rect -25 305 -5 375
rect 115 620 135 690
rect 220 620 240 690
<< psubdiff >>
rect 140 -130 240 -115
rect 140 -150 155 -130
rect 225 -150 240 -130
rect 140 -165 240 -150
<< nsubdiff >>
rect 20 860 70 875
rect 20 790 35 860
rect 55 790 70 860
rect 20 775 70 790
<< psubdiffcont >>
rect 155 -150 225 -130
<< nsubdiffcont >>
rect 35 790 55 860
<< poly >>
rect -75 875 -60 890
rect 150 875 165 890
rect 190 875 205 890
rect -75 765 -60 775
rect -75 750 90 765
rect -55 705 -40 720
rect -55 575 -40 605
rect -55 560 35 575
rect -55 520 -40 535
rect -55 390 -40 420
rect -55 235 -40 290
rect 20 260 35 560
rect -5 245 35 260
rect -5 235 10 245
rect -5 120 10 135
rect -5 110 40 120
rect -5 90 10 110
rect 30 90 40 110
rect -5 80 40 90
rect 75 55 90 750
rect 150 705 165 775
rect 190 760 205 775
rect 190 750 280 760
rect 190 745 250 750
rect 240 730 250 745
rect 270 730 280 750
rect 240 720 280 730
rect 190 705 205 720
rect 150 520 165 605
rect 190 575 205 605
rect 190 565 240 575
rect 190 545 200 565
rect 220 545 240 565
rect 190 535 240 545
rect 150 390 165 420
rect 150 240 165 290
rect 225 240 240 535
rect -5 45 90 55
rect -5 25 5 45
rect 25 40 90 45
rect 115 225 165 240
rect 190 225 240 240
rect 25 25 35 40
rect -5 15 35 25
rect -5 -65 10 15
rect -55 -190 -40 -165
rect -5 -180 10 -165
rect 115 -190 130 225
rect 190 215 205 225
rect 190 100 205 115
rect 190 90 230 100
rect 190 70 200 90
rect 220 70 230 90
rect 190 60 230 70
rect 190 20 205 35
rect 190 -90 205 -80
rect 265 -90 280 720
rect 190 -105 280 -90
rect -80 -200 -40 -190
rect -80 -220 -70 -200
rect -50 -220 -40 -200
rect -80 -230 -40 -220
rect 90 -200 130 -190
rect 90 -220 100 -200
rect 120 -220 130 -200
rect 90 -230 130 -220
<< polycont >>
rect 10 90 30 110
rect 250 730 270 750
rect 200 545 220 565
rect 5 25 25 45
rect 200 70 220 90
rect -70 -220 -50 -200
rect 100 -220 120 -200
<< locali >>
rect -120 860 -80 870
rect -120 790 -110 860
rect -90 790 -80 860
rect -120 780 -80 790
rect -55 860 -15 870
rect -55 790 -45 860
rect -25 790 -15 860
rect -55 780 -15 790
rect 25 860 65 870
rect 25 790 35 860
rect 55 800 65 860
rect 105 860 145 870
rect 105 800 115 860
rect 55 790 115 800
rect 135 790 145 860
rect 210 860 250 870
rect 210 800 220 860
rect 25 780 145 790
rect -100 700 -80 780
rect -35 760 -15 780
rect -35 740 85 760
rect -100 690 -60 700
rect -100 620 -90 690
rect -70 620 -60 690
rect -100 610 -60 620
rect -35 690 5 700
rect -35 620 -25 690
rect -5 630 5 690
rect -5 620 45 630
rect -35 610 45 620
rect -100 505 -60 515
rect -100 435 -90 505
rect -70 435 -60 505
rect -100 425 -60 435
rect -35 505 5 515
rect -35 435 -25 505
rect -5 435 5 505
rect -35 425 5 435
rect 25 385 45 610
rect -100 375 -60 385
rect -100 305 -90 375
rect -70 305 -60 375
rect -100 295 -60 305
rect -35 375 45 385
rect -35 305 -25 375
rect -5 365 45 375
rect -5 305 5 365
rect -35 295 5 305
rect 25 230 45 365
rect 65 445 85 740
rect 125 700 145 780
rect 105 690 145 700
rect 105 620 115 690
rect 135 620 145 690
rect 105 610 145 620
rect 170 790 220 800
rect 240 790 250 860
rect 170 780 250 790
rect 170 575 190 780
rect 240 750 280 760
rect 240 740 250 750
rect 220 730 250 740
rect 270 730 280 750
rect 220 720 280 730
rect 220 700 240 720
rect 210 690 250 700
rect 210 620 220 690
rect 240 630 250 690
rect 240 620 270 630
rect 210 610 270 620
rect 170 565 230 575
rect 170 545 200 565
rect 220 545 230 565
rect 170 535 230 545
rect 170 515 190 535
rect 105 505 145 515
rect 105 445 115 505
rect 65 435 115 445
rect 135 435 145 505
rect 65 425 145 435
rect 170 505 210 515
rect 170 435 180 505
rect 200 435 210 505
rect 170 425 210 435
rect 65 270 85 425
rect 105 375 145 385
rect 105 305 115 375
rect 135 305 145 375
rect 105 295 145 305
rect 170 375 210 385
rect 170 305 180 375
rect 200 315 210 375
rect 250 315 270 610
rect 200 305 270 315
rect 170 295 270 305
rect 65 250 95 270
rect -100 220 -60 230
rect -100 -150 -90 220
rect -70 -150 -60 220
rect 15 220 55 230
rect 15 160 25 220
rect -40 150 25 160
rect 45 150 55 220
rect -40 140 55 150
rect -40 55 -20 140
rect 75 120 95 250
rect 250 210 270 295
rect 145 200 185 210
rect 145 130 155 200
rect 175 130 185 200
rect 145 120 185 130
rect 210 200 270 210
rect 210 130 220 200
rect 240 190 270 200
rect 240 130 250 190
rect 210 120 250 130
rect 0 110 95 120
rect 0 90 10 110
rect 30 100 95 110
rect 30 90 40 100
rect 0 80 40 90
rect -40 45 35 55
rect -40 35 5 45
rect -5 25 5 35
rect 25 25 35 45
rect -5 15 35 25
rect 75 -70 95 100
rect 190 90 230 100
rect 190 70 200 90
rect 220 70 230 90
rect 190 60 230 70
rect 210 15 230 60
rect -100 -160 -60 -150
rect 15 -80 95 -70
rect 15 -150 25 -80
rect 45 -90 95 -80
rect 145 5 185 15
rect 145 -65 155 5
rect 175 -65 185 5
rect 145 -75 185 -65
rect 210 5 250 15
rect 210 -65 220 5
rect 240 -65 250 5
rect 210 -75 250 -65
rect 45 -150 55 -90
rect 15 -160 55 -150
rect 145 -120 165 -75
rect 145 -130 235 -120
rect 145 -150 155 -130
rect 225 -150 235 -130
rect 145 -160 235 -150
rect -80 -200 -40 -190
rect -80 -220 -70 -200
rect -50 -220 -40 -200
rect -80 -230 -40 -220
rect 90 -200 130 -190
rect 90 -220 100 -200
rect 120 -220 130 -200
rect 90 -230 130 -220
<< viali >>
rect -110 790 -90 860
rect 35 790 55 860
rect 115 790 135 860
rect -90 620 -70 690
rect -90 435 -70 505
rect -25 435 -5 505
rect -90 305 -70 375
rect -25 305 -5 375
rect 115 620 135 690
rect 115 435 135 505
rect 180 435 200 505
rect 115 305 135 375
rect 180 305 200 375
rect -90 -150 -70 220
rect 155 130 175 200
rect 155 -65 175 5
rect 155 -150 225 -130
rect -70 -220 -50 -200
rect 100 -220 120 -200
<< metal1 >>
rect -125 860 280 895
rect -125 790 -110 860
rect -90 790 35 860
rect 55 790 115 860
rect 135 790 280 860
rect -125 690 280 790
rect -125 620 -90 690
rect -70 620 115 690
rect 135 620 280 690
rect -125 585 280 620
rect -125 505 -60 520
rect -125 435 -90 505
rect -70 435 -60 505
rect -125 420 -60 435
rect -35 505 145 520
rect -35 435 -25 505
rect -5 435 115 505
rect 135 435 145 505
rect -35 420 145 435
rect 170 505 280 520
rect 170 435 180 505
rect 200 435 280 505
rect 170 420 280 435
rect -125 375 -60 390
rect -125 305 -90 375
rect -70 305 -60 375
rect -125 290 -60 305
rect -35 375 145 390
rect -35 305 -25 375
rect -5 305 115 375
rect 135 305 145 375
rect -35 290 145 305
rect 170 375 280 390
rect 170 305 180 375
rect 200 305 280 375
rect 170 290 280 305
rect -125 220 280 235
rect -125 -150 -90 220
rect -70 200 280 220
rect -70 130 155 200
rect 175 130 280 200
rect -70 5 280 130
rect -70 -65 155 5
rect 175 -65 280 5
rect -70 -130 280 -65
rect -70 -150 155 -130
rect 225 -150 280 -130
rect -125 -160 280 -150
rect -125 -200 280 -190
rect -125 -220 -70 -200
rect -50 -220 100 -200
rect 120 -220 280 -200
rect -125 -230 280 -220
<< labels >>
rlabel metal1 -125 -210 -125 -210 7 CLK
port 1 w
rlabel metal1 -125 35 -125 35 7 VN
port 2 w
rlabel metal1 -125 340 -125 340 7 Dn
port 3 w
rlabel metal1 -125 470 -125 470 7 D
port 4 w
rlabel metal1 -125 735 -125 735 7 VP
port 5 w
rlabel metal1 280 470 280 470 3 Q
port 6 e
rlabel metal1 280 340 280 340 3 Qn
port 7 e
<< end >>
